// PE_tb.v
// Testbench for PE


module PE_tb();

    

endmodule