// PEarray.v
//  systolic array 

module PEarray#(
    parameter DATA_WIDTH = 8,
    parameter PE_CHANNEL = 4,
    parameter PE_ROW = 25
)(
    input clk,
    input rst_n,
    input mode
);




endmodule