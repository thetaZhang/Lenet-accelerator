// InputDataBuffer.v
// Input data buffer, reorder with the shape of conv kernel

module InputDataBuffer#(
    parameter DATA_WIDTH = 8,
    parameter 
)(

);



endmodule